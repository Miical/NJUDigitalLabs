module bcd7seg(
  input [3:0] b,
  input en,
  output reg [7:0] h
);

  always @(*) begin
    if (!en) begin
      h = 8'b11111111;
    end else case(b)
      4'b0000: h = 8'b11000000;
      4'b0001: h = 8'b11111001;
      4'b0010: h = 8'b10100100;
      4'b0011: h = 8'b10110000;
      4'b0100: h = 8'b10011001;
      4'b0101: h = 8'b10010010;
      4'b0110: h = 8'b10000010;
      4'b0111: h = 8'b11111000;
      4'b1000: h = 8'b10000000;
      4'b1001: h = 8'b10010000;
      4'b1010: h = 8'b10001000;
      4'b1011: h = 8'b10000011;
      4'b1100: h = 8'b11000110;
      4'b1101: h = 8'b10100001;
      4'b1110: h = 8'b10000110;
      4'b1111: h = 8'b10001110;
      default: h = 8'b11111111;
    endcase
  end

endmodule
